module dffer(D,clk,E,R,Q);
input D;      // Data input 
input clk;    // clock input 
input E;      // enable 
input R;      // reset input 
output Q;     // output Q 

endmodule 
