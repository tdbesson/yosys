module dffe(D,clk,E,Q);
input D;     // Data input 
input clk;   // clock input 
input E;     //  enable
output Q;    // output Q 

endmodule 
