module dffes(D,clk,E,S,Q);
input D;      // Data input 
input clk;    // clock input 
input E;      // enable 
input S;      // set input 
output Q;     // output Q 

endmodule 
