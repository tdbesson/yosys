module dffs(D,clk,S,Q);
input D;      // Data input 
input clk;    // clock input 
input S;      // set input 
output Q;     // output Q 

endmodule 
