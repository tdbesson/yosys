module dffers(D,clk,E,R,S,Q);
input D;      // Data input 
input clk;    // clock input 
input E;      // enable 
input R;      // reset input 
input S;      // set input 
output Q;     // output Q 

endmodule 
