module dffrs(D,clk,R,S,Q);
input D;      // Data input 
input clk;    // clock input 
input R;      // reset input 
input S;      // set input 
output Q;     // output Q 

endmodule 
