module dffr(D,clk,R,Q);
input D;      // Data input 
input clk;    // clock input 
input R;      // reset input 
output Q;     // output Q 

endmodule 
